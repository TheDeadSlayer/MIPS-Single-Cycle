`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:13:00 06/03/2021 
// Design Name: 
// Module Name:    PC_MahmoudSaeed_18102867 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module PC_MahmoudSaeed_18102867(
    input [31:0] PCin,
    input CLK,
    input [31:0] PCout
    );


endmodule
